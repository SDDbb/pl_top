`timescale 1ns/1ps

// =====================================================================
// btn_start_gen
// ʹ�ð��ذ�������"��ʼһ֡"�ĵ��������� start_pulse
//
// ���ܣ�
// 1) ���첽��������ͬ���� clk ��
// 2) �� 10ms ȥ�������õ��ȶ�������ƽ btn_stable
// 3) �� btn_stable ������������⣬��� 1clk ��ȵ� start_pulse
//
// ˵����
// - ���谴��Ϊ����Ч������ = 0���ɿ� = 1
//   �����İ����Ǹ���Ч���� button_level = ~button_sync2 �ĳ� button_level = button_sync2
// =====================================================================
module btn_start_gen #(
    parameter integer CLK_FREQ_HZ     = 50_000_000, // ʱ��Ƶ��
    parameter integer DEBOUNCE_MS     = 10          // ȥ��ʱ�� (ms)
)(
    input  wire clk,
    input  wire rst_n,         // ����Ч��λ

    input  wire button_in,     // ���� PL ������ԭʼ�ź�
    output wire start_pulse    // 1 �� clk ���ڵ���������
);

    // --------------------------------------------------------------
    // 1. ����ͬ���� clk ��
    // --------------------------------------------------------------
    reg button_sync1, button_sync2;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            button_sync1 <= 1'b1;
            button_sync2 <= 1'b1;
        end else begin
            button_sync1 <= button_in;
            button_sync2 <= button_sync1;
        end
    end

    // ���谴��Ϊ����Ч������=0���ɿ�=1
    // ������Ч���ĳ� button_level = button_sync2;
    wire button_level = ~button_sync2;

    // --------------------------------------------------------------
    // 2. ȥ����ֻ�е���ƽ�����ȶ� DEBOUNCE_MS ����Ϊ״̬�ı�
    // --------------------------------------------------------------
    localparam integer DEBOUNCE_CNT_MAX =
        (CLK_FREQ_HZ / 1000) * DEBOUNCE_MS;

    localparam integer DEBOUNCE_CNT_BITS =
        $clog2(DEBOUNCE_CNT_MAX+1);

    reg [DEBOUNCE_CNT_BITS-1:0] db_cnt;
    reg                         btn_stable;      // ȥ������ȶ�������ƽ

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            db_cnt    <= {DEBOUNCE_CNT_BITS{1'b0}};
            btn_stable <= 1'b0;
        end else begin
            // �����ǰ�����İ�����ƽ����һ���ȶ�ֵ��ͬ �� ���¼�ʱ
            if (button_level != btn_stable) begin
                if (db_cnt < DEBOUNCE_CNT_MAX[DEBOUNCE_CNT_BITS-1:0]) begin
                    db_cnt <= db_cnt + 1'b1;
                end else begin
                    // ��ƽ�Ѿ��ȶ�����ȥ��ʱ�� �� �����ȶ�ֵ
                    btn_stable <= button_level;
                    db_cnt     <= {DEBOUNCE_CNT_BITS{1'b0}};
                end
            end else begin
                // ��ƽû�䣬��������
                db_cnt <= {DEBOUNCE_CNT_BITS{1'b0}};
            end
        end
    end

    // --------------------------------------------------------------
    // 3. �����ؼ�⣺��"δ����"��"����"��˲����� 1clk ����
    //    ��ÿ��һ�μ�ֻ����һ�� start_pulse��
    // --------------------------------------------------------------
    reg btn_stable_d;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            btn_stable_d <= 1'b0;
        else
            btn_stable_d <= btn_stable;
    end

    assign start_pulse = btn_stable & ~btn_stable_d;

endmodule
