`timescale 1ns/1ps

// -----------------------------------------------------------------------------
// rx_photon_frontend (improved robust version)
// -----------------------------------------------------------------------------
// ���ܣ�
// 1) �����ԱȽ������첽 SPAD ����ͬ���� clk_sys
// 2) ���� 1clk ��ȵ� photon event pulse
//
// �Ľ��㣨�����ԭ�棩��
// - USE_HOLDOFF=0 ʱ����ȫ��ȥ�أ�spad_pulse_sync = raw_evt��
// - HOLD_CYCLES=0 ʱ����ʹ USE_HOLDOFF=1��Ҳ����ǿ�Ʋ��� 1clk ����
//   ��HOLD=0 ����"������"��
// -----------------------------------------------------------------------------

module rx_photon_frontend (
    input  wire clk_sys,          // ϵͳʱ�ӣ��� 130 MHz��
    input  wire rst_n,

    input  wire spad_pulse_in,     // ���ԱȽ������첽��������
    output wire spad_pulse_sync    // ͬ����� 1clk ���壨�����¼���
);

    // ------------------------------------------------------------
    // 1) ˫������ͬ����CDC��
    // ------------------------------------------------------------
    (* ASYNC_REG = "TRUE" *) reg spad_ff1;
    (* ASYNC_REG = "TRUE" *) reg spad_ff2;

    always @(posedge clk_sys or negedge rst_n) begin
        if (!rst_n) begin
            spad_ff1 <= 1'b0;
            spad_ff2 <= 1'b0;
        end else begin
            spad_ff1 <= spad_pulse_in;
            spad_ff2 <= spad_ff1;
        end
    end
    
    assign spad_pulse_sync = spad_ff2;
endmodule
