`timescale 1ns/1ps

// ============================================================
// cdc_pulse_sync
// ���ܣ�
//   �� src_clk ��� 1clk ���壬��ȫ��ͬ���� dst_clk ��
//   ���� dst_clk ����� 1clk ��ȵ�����
//
// ԭ��
//   - Դ�򣺰� pulse ��ת�� toggle
//   - Ŀ���򣺶� toggle ������
//   - ��� toggle ��ת �� ���� 1clk pulse
// ============================================================
module cdc_pulse_sync (
    input  wire src_clk,
    input  wire src_rst_n,
    input  wire src_pulse,   // src_clk ��� 1clk ����

    input  wire dst_clk,
    input  wire dst_rst_n,
    output wire dst_pulse    // dst_clk ��� 1clk ����
);

    // ------------------------------------------------
    // Դʱ����pulse �� toggle
    // ------------------------------------------------
    reg src_toggle;

    always @(posedge src_clk or negedge src_rst_n) begin
        if (!src_rst_n)
            src_toggle <= 1'b0;
        else if (src_pulse)
            src_toggle <= ~src_toggle;
    end

    // ------------------------------------------------
    // Ŀ��ʱ����ͬ�� toggle
    // ------------------------------------------------
    reg dst_toggle_ff1, dst_toggle_ff2;

    always @(posedge dst_clk or negedge dst_rst_n) begin
        if (!dst_rst_n) begin
            dst_toggle_ff1 <= 1'b0;
            dst_toggle_ff2 <= 1'b0;
        end else begin
            dst_toggle_ff1 <= src_toggle;
            dst_toggle_ff2 <= dst_toggle_ff1;
        end
    end

    // ------------------------------------------------
    // toggle ���ؼ�� �� 1clk pulse
    // ------------------------------------------------
    assign dst_pulse = dst_toggle_ff1 ^ dst_toggle_ff2;

endmodule
